 module time_stamp
 (
 output wire [31:0]  time_dout
);
 assign time_dout  = 32'd1513122301;
 endmodule
